package States;
typedef enum logic [3:0] { EXACT, OVERFLOW, UNDERFLOW, INEXACT } State_e;
endpackage
